module alu_ov (a,b,aluc,r,z,v); // 32-bit alu with zero and overflow flags
input [31:0] a, b; // inputs: a, b
input [3:0] aluc; // input: alu control: // aluc[3:0]:
output [31:0] r; // output: alu result // x 0 0 0 ADD
output z, v; // outputs: zero, overflow // x 1 0 0 SUB
wire [31:0] d_and = a & b; // x 0 0 1 AND
wire [31:0] d_or = a | b; // x 1 0 1 OR
wire [31:0] d_xor = a ^ b; // x 0 1 0 XOR
wire [31:0] d_lui = {b[15:0],16'h0}; // x 1 1 0 LUI
wire [31:0] d_and_or = aluc[2]? d_or : d_and; // 0 0 1 1 SLL
wire [31:0] d_xor_lui = aluc[2]? d_lui : d_xor; // 0 1 1 1 SRL
wire [31:0] d_as,d_sh; // 1 1 1 1 SRA
// addsub32 (a,b,sub, s);
addsub32 as32 (a,b,aluc[2],d_as); // add/sub
// shift (d,sa, right, arith, sh);
shift shifter (b,a[4:0],aluc[2],aluc[3],d_sh); // shift
// mux4x32 (a0, a1, a2, a3, s, y);
mux4x32 res (d_as,d_and_or,d_xor_lui,d_sh,aluc[1:0],r); // alu result
assign z = ~|r; // z = (r == 0)
assign v = ~aluc[2] & ~a[31] & ~b[31] & r[31] & ~aluc[1] & ~aluc[0] | ~aluc[2] & a[31] & b[31] & ~r[31] & ~aluc[1] & ~aluc[0] | aluc[2] & ~a[31] & b[31] & r[31] & ~aluc[1] & ~aluc[0] | aluc[2] & a[31] & ~b[31] & ~r[31] & ~aluc[1] & ~aluc[0];
endmodule